module cosineTable (
    input [7:0] angle,             // 8-bit angle input (0-255, 0 to 360 degrees)
    output reg signed [15:0] cosine  // 16-bit signed output value (scaled by 8192)
);

always @(*) begin
    case(angle)
        8'h00: cosine = 16'h3fff ;
        8'h01: cosine = 16'h3ffa ;
        8'h02: cosine = 16'h3feb ;
        8'h03: cosine = 16'h3fd2 ;
        8'h04: cosine = 16'h3fb0 ;
        8'h05: cosine = 16'h3f83 ;
        8'h06: cosine = 16'h3f4d ;
        8'h07: cosine = 16'h3f0d ;
        8'h08: cosine = 16'h3ec4 ;
        8'h09: cosine = 16'h3e70 ;
        8'h0a: cosine = 16'h3e14 ;
        8'h0b: cosine = 16'h3dad ;
        8'h0c: cosine = 16'h3d3d ;
        8'h0d: cosine = 16'h3cc4 ;
        8'h0e: cosine = 16'h3c41 ;
        8'h0f: cosine = 16'h3bb5 ;
        8'h10: cosine = 16'h3b1f ;
        8'h11: cosine = 16'h3a81 ;
        8'h12: cosine = 16'h39da ;
        8'h13: cosine = 16'h3929 ;
        8'h14: cosine = 16'h3870 ;
        8'h15: cosine = 16'h37ae ;
        8'h16: cosine = 16'h36e4 ;
        8'h17: cosine = 16'h3611 ;
        8'h18: cosine = 16'h3535 ;
        8'h19: cosine = 16'h3452 ;
        8'h1a: cosine = 16'h3366 ;
        8'h1b: cosine = 16'h3273 ;
        8'h1c: cosine = 16'h3178 ;
        8'h1d: cosine = 16'h3075 ;
        8'h1e: cosine = 16'h2f6b ;
        8'h1f: cosine = 16'h2e59 ;
        8'h20: cosine = 16'h2d40 ;
        8'h21: cosine = 16'h2c20 ;
        8'h22: cosine = 16'h2afa ;
        8'h23: cosine = 16'h29cc ;
        8'h24: cosine = 16'h2899 ;
        8'h25: cosine = 16'h275f ;
        8'h26: cosine = 16'h261f ;
        8'h27: cosine = 16'h24d9 ;
        8'h28: cosine = 16'h238d ;
        8'h29: cosine = 16'h223c ;
        8'h2a: cosine = 16'h20e6 ;
        8'h2b: cosine = 16'h1f8b ;
        8'h2c: cosine = 16'h1e2a ;
        8'h2d: cosine = 16'h1cc5 ;
        8'h2e: cosine = 16'h1b5c ;
        8'h2f: cosine = 16'h19ef ;
        8'h30: cosine = 16'h187d ;
        8'h31: cosine = 16'h1708 ;
        8'h32: cosine = 16'h158f ;
        8'h33: cosine = 16'h1413 ;
        8'h34: cosine = 16'h1293 ;
        8'h35: cosine = 16'h1111 ;
        8'h36: cosine = 16'h0f8c ;
        8'h37: cosine = 16'h0e05 ;
        8'h38: cosine = 16'h0c7c ;
        8'h39: cosine = 16'h0af0 ;
        8'h3a: cosine = 16'h0963 ;
        8'h3b: cosine = 16'h07d5 ;
        8'h3c: cosine = 16'h0645 ;
        8'h3d: cosine = 16'h04b5 ;
        8'h3e: cosine = 16'h0323 ;
        8'h3f: cosine = 16'h0192 ;
        8'h40: cosine = 16'h0000 ;
        8'h41: cosine = 16'hfe6e ;
        8'h42: cosine = 16'hfcdd ;
        8'h43: cosine = 16'hfb4b ;
        8'h44: cosine = 16'hf9bb ;
        8'h45: cosine = 16'hf82b ;
        8'h46: cosine = 16'hf69d ;
        8'h47: cosine = 16'hf510 ;
        8'h48: cosine = 16'hf384 ;
        8'h49: cosine = 16'hf1fb ;
        8'h4a: cosine = 16'hf074 ;
        8'h4b: cosine = 16'heeef ;
        8'h4c: cosine = 16'hed6d ;
        8'h4d: cosine = 16'hebed ;
        8'h4e: cosine = 16'hea71 ;
        8'h4f: cosine = 16'he8f8 ;
        8'h50: cosine = 16'he783 ;
        8'h51: cosine = 16'he611 ;
        8'h52: cosine = 16'he4a4 ;
        8'h53: cosine = 16'he33b ;
        8'h54: cosine = 16'he1d6 ;
        8'h55: cosine = 16'he075 ;
        8'h56: cosine = 16'hdf1a ;
        8'h57: cosine = 16'hddc4 ;
        8'h58: cosine = 16'hdc73 ;
        8'h59: cosine = 16'hdb27 ;
        8'h5a: cosine = 16'hd9e1 ;
        8'h5b: cosine = 16'hd8a1 ;
        8'h5c: cosine = 16'hd767 ;
        8'h5d: cosine = 16'hd634 ;
        8'h5e: cosine = 16'hd506 ;
        8'h5f: cosine = 16'hd3e0 ;
        8'h60: cosine = 16'hd2c0 ;
        8'h61: cosine = 16'hd1a7 ;
        8'h62: cosine = 16'hd095 ;
        8'h63: cosine = 16'hcf8b ;
        8'h64: cosine = 16'hce88 ;
        8'h65: cosine = 16'hcd8d ;
        8'h66: cosine = 16'hcc9a ;
        8'h67: cosine = 16'hcbae ;
        8'h68: cosine = 16'hcacb ;
        8'h69: cosine = 16'hc9ef ;
        8'h6a: cosine = 16'hc91c ;
        8'h6b: cosine = 16'hc852 ;
        8'h6c: cosine = 16'hc790 ;
        8'h6d: cosine = 16'hc6d7 ;
        8'h6e: cosine = 16'hc626 ;
        8'h6f: cosine = 16'hc57f ;
        8'h70: cosine = 16'hc4e1 ;
        8'h71: cosine = 16'hc44b ;
        8'h72: cosine = 16'hc3bf ;
        8'h73: cosine = 16'hc33c ;
        8'h74: cosine = 16'hc2c3 ;
        8'h75: cosine = 16'hc253 ;
        8'h76: cosine = 16'hc1ec ;
        8'h77: cosine = 16'hc190 ;
        8'h78: cosine = 16'hc13c ;
        8'h79: cosine = 16'hc0f3 ;
        8'h7a: cosine = 16'hc0b3 ;
        8'h7b: cosine = 16'hc07d ;
        8'h7c: cosine = 16'hc050 ;
        8'h7d: cosine = 16'hc02e ;
        8'h7e: cosine = 16'hc015 ;
        8'h7f: cosine = 16'hc006 ;
        8'h80: cosine = 16'hc001 ;
        8'h81: cosine = 16'hc006 ;
        8'h82: cosine = 16'hc015 ;
        8'h83: cosine = 16'hc02e ;
        8'h84: cosine = 16'hc050 ;
        8'h85: cosine = 16'hc07d ;
        8'h86: cosine = 16'hc0b3 ;
        8'h87: cosine = 16'hc0f3 ;
        8'h88: cosine = 16'hc13c ;
        8'h89: cosine = 16'hc190 ;
        8'h8a: cosine = 16'hc1ec ;
        8'h8b: cosine = 16'hc253 ;
        8'h8c: cosine = 16'hc2c3 ;
        8'h8d: cosine = 16'hc33c ;
        8'h8e: cosine = 16'hc3bf ;
        8'h8f: cosine = 16'hc44b ;
        8'h90: cosine = 16'hc4e1 ;
        8'h91: cosine = 16'hc57f ;
        8'h92: cosine = 16'hc626 ;
        8'h93: cosine = 16'hc6d7 ;
        8'h94: cosine = 16'hc790 ;
        8'h95: cosine = 16'hc852 ;
        8'h96: cosine = 16'hc91c ;
        8'h97: cosine = 16'hc9ef ;
        8'h98: cosine = 16'hcacb ;
        8'h99: cosine = 16'hcbae ;
        8'h9a: cosine = 16'hcc9a ;
        8'h9b: cosine = 16'hcd8d ;
        8'h9c: cosine = 16'hce88 ;
        8'h9d: cosine = 16'hcf8b ;
        8'h9e: cosine = 16'hd095 ;
        8'h9f: cosine = 16'hd1a7 ;
        8'ha0: cosine = 16'hd2c0 ;
        8'ha1: cosine = 16'hd3e0 ;
        8'ha2: cosine = 16'hd506 ;
        8'ha3: cosine = 16'hd634 ;
        8'ha4: cosine = 16'hd767 ;
        8'ha5: cosine = 16'hd8a1 ;
        8'ha6: cosine = 16'hd9e1 ;
        8'ha7: cosine = 16'hdb27 ;
        8'ha8: cosine = 16'hdc73 ;
        8'ha9: cosine = 16'hddc4 ;
        8'haa: cosine = 16'hdf1a ;
        8'hab: cosine = 16'he075 ;
        8'hac: cosine = 16'he1d6 ;
        8'had: cosine = 16'he33b ;
        8'hae: cosine = 16'he4a4 ;
        8'haf: cosine = 16'he611 ;
        8'hb0: cosine = 16'he783 ;
        8'hb1: cosine = 16'he8f8 ;
        8'hb2: cosine = 16'hea71 ;
        8'hb3: cosine = 16'hebed ;
        8'hb4: cosine = 16'hed6d ;
        8'hb5: cosine = 16'heeef ;
        8'hb6: cosine = 16'hf074 ;
        8'hb7: cosine = 16'hf1fb ;
        8'hb8: cosine = 16'hf384 ;
        8'hb9: cosine = 16'hf510 ;
        8'hba: cosine = 16'hf69d ;
        8'hbb: cosine = 16'hf82b ;
        8'hbc: cosine = 16'hf9bb ;
        8'hbd: cosine = 16'hfb4b ;
        8'hbe: cosine = 16'hfcdd ;
        8'hbf: cosine = 16'hfe6e ;
        8'hc0: cosine = 16'h0000 ;
        8'hc1: cosine = 16'h0192 ;
        8'hc2: cosine = 16'h0323 ;
        8'hc3: cosine = 16'h04b5 ;
        8'hc4: cosine = 16'h0645 ;
        8'hc5: cosine = 16'h07d5 ;
        8'hc6: cosine = 16'h0963 ;
        8'hc7: cosine = 16'h0af0 ;
        8'hc8: cosine = 16'h0c7c ;
        8'hc9: cosine = 16'h0e05 ;
        8'hca: cosine = 16'h0f8c ;
        8'hcb: cosine = 16'h1111 ;
        8'hcc: cosine = 16'h1293 ;
        8'hcd: cosine = 16'h1413 ;
        8'hce: cosine = 16'h158f ;
        8'hcf: cosine = 16'h1708 ;
        8'hd0: cosine = 16'h187d ;
        8'hd1: cosine = 16'h19ef ;
        8'hd2: cosine = 16'h1b5c ;
        8'hd3: cosine = 16'h1cc5 ;
        8'hd4: cosine = 16'h1e2a ;
        8'hd5: cosine = 16'h1f8b ;
        8'hd6: cosine = 16'h20e6 ;
        8'hd7: cosine = 16'h223c ;
        8'hd8: cosine = 16'h238d ;
        8'hd9: cosine = 16'h24d9 ;
        8'hda: cosine = 16'h261f ;
        8'hdb: cosine = 16'h275f ;
        8'hdc: cosine = 16'h2899 ;
        8'hdd: cosine = 16'h29cc ;
        8'hde: cosine = 16'h2afa ;
        8'hdf: cosine = 16'h2c20 ;
        8'he0: cosine = 16'h2d40 ;
        8'he1: cosine = 16'h2e59 ;
        8'he2: cosine = 16'h2f6b ;
        8'he3: cosine = 16'h3075 ;
        8'he4: cosine = 16'h3178 ;
        8'he5: cosine = 16'h3273 ;
        8'he6: cosine = 16'h3366 ;
        8'he7: cosine = 16'h3452 ;
        8'he8: cosine = 16'h3535 ;
        8'he9: cosine = 16'h3611 ;
        8'hea: cosine = 16'h36e4 ;
        8'heb: cosine = 16'h37ae ;
        8'hec: cosine = 16'h3870 ;
        8'hed: cosine = 16'h3929 ;
        8'hee: cosine = 16'h39da ;
        8'hef: cosine = 16'h3a81 ;
        8'hf0: cosine = 16'h3b1f ;
        8'hf1: cosine = 16'h3bb5 ;
        8'hf2: cosine = 16'h3c41 ;
        8'hf3: cosine = 16'h3cc4 ;
        8'hf4: cosine = 16'h3d3d ;
        8'hf5: cosine = 16'h3dad ;
        8'hf6: cosine = 16'h3e14 ;
        8'hf7: cosine = 16'h3e70 ;
        8'hf8: cosine = 16'h3ec4 ;
        8'hf9: cosine = 16'h3f0d ;
        8'hfa: cosine = 16'h3f4d ;
        8'hfb: cosine = 16'h3f83 ;
        8'hfc: cosine = 16'h3fb0 ;
        8'hfd: cosine = 16'h3fd2 ;
        8'hfe: cosine = 16'h3feb ;
        8'hff: cosine = 16'h3ffa ;
    endcase
end
   
endmodule
